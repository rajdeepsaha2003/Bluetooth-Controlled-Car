PK   ���W��1W  �    cirkitFile.json�]�7��W�W���c�%�]\�����؆��Xر��h�d��G������*J���Xdg��b5�c�����ا���u�ۗ�_���f�]<P�\�K�����d���ٮ�����û��'�{r��C���v�r{X��X+�NRY��P$K�eb��rͤ�Ԯ��������)�;�u���u�
�2Q�6Os?eF��ʍPEFi����#��ȂXn���̍L�M,Qi����*���P�d�Wy�R��D�p�"1:IaE�!�h�fl�/��p�,W��$M�ȍ�kܸD���YF2�ʤ�1[*0[�rU)�����,��P:a�Ȣ�&Í�#��Z`F68h[�ƪ�^�H�@���
d�쯐�C�M�͵Ty�˜$�0<I�	%���Dr䖡H�R������b�f��Y`h�b�M8�hv��!�R�7v����ƭvȘ��ƁeN)ʞ2�[���4��
36GZr�� �C*��"'���,s�Q���y��,�J��S��yÌ2���C
�-h^�D�~B����I��gy�)fq�ҧ��1rH��l��!e��L�b)�37��*Kܙ��4�EU�l�T)hd�4nS�]4P�ppۘa�5�����_�ب-FQ������b�Fmp��PÏ;�ǡ�xl�W�&�B��&�#�9�d`�:��AC�S���L70���FA�(����!��!b�P�9�S�Ę f8w�*7�ڰ������s�,+TR�DZ2��*���!u ��:�s��ZK�VZ�����&B*���"!i�����yp���4B���H��\�^<P�D.�-u���-n� f�f����Y*uQ��B��([$��HBJ�ӔɼJ���3��-B��lÞ�@�op~@�0Bk��*���I&+�Xj�)�<%y|f�	)h��3�R�@��GN�!uh����:l	xp��l�.����L\�o?������yee���!V�F�¢p�Q��%�H.2�,*
�TU)	Cp1Qd�qP	�q�K�����/q��A0�aZc�*���&��=�(-��M0�E��W���g6�(a����#�*�Ql*�L�؜P��,҂�8�P����9��J!0lN��r]b��(���b؜t��x ���0ޓ�zPDr�#�䆂FG�EL� �C��ԛ)-�\tY&�(7�i�|�;�:�g��|�:�:�'��|:�:���z49�����z�8�D@�=�`�y�TV�c�\�)��E�G�ɘz��2��Ӣq�=�"�iʸ,Г�qY���L���a<���o����,�<��,М��A�������[��R�T�,д�9�}��>�C���n���>}Df`�\X.<
����EEᢣp1Q��8���8�q�K����0��`�4�i�8(fqP�"��8(fqP�⠘�A1��b�,�Y�8(�(g`�\��2���X<������Ln&p�er+�3�P	�q�;���3����W����g`�\&����s�\lp�er��X<��5g`�\��2�p�e��X<�IY�X<�IY�X<�i-���L����L����L����Lk)h��R��K�㯇�����u���r�q�/��Ӽ,֛�z�/����u�7���Uc�1�J`d������@����##3Lf��,p{ �FTE7ʋG�����U����Pc#/��F]�����.&�wO�#��G��6�4z}2�2z�1�Sǉq�1#c����Lx`Nwo���g���0�t#�BC�5�!fhd����)G�op�q�zLp�+�fvcFFנFh�"��c�P�K`n��`�����&��/��~)�u�-�r���_,����y�Q�~�Y�Q�c ��� 65Al�"��DE���"`��"�#{� �ĸ� �\�͖ ����edf/ 2�1*�=�x��Q����{��3�́�%��B�%�GF/61r3	����-4M2*�=�%��#i� �;��DQ�wɤ���wH��\����2s������"�ϛ��������}������1�ٟ!�sd����QL�C�ء_��f�0�M���8.9��=4x��X�R,~���(�@a�aI�oSC	d��n�r��@^���z��üz����-�K�:z%߀�� ���4A�e@O��b��Px���1�����v6@�0��;�0�7�oO������
�7����&žԭ��7�H���&p=!�����!�,7�dn ܨc�t#�̠�^g��:��=]�<�\s��oq<L����#.G�L<ZW$Fd7��q� ���.`�U����+v. �p��.`T��v���2v�a�*�\��\�[Yp�#le�u�v�W�u�ᾍ�Z	�\I:���xF�jI�t�I�t���6�Pf\H�aW���ͦ��n��ɧ�!a�����1/�߱~�y_�;��{�x4�i�5D�u��]o��q�ݍ�I��V÷��:�Q?3�=�3��RP}9��$U_֪/�՗׸�����@\������G�1�8/\��m��:A�ck��ju��V�^ou���v��ku�(�V��h/`�^tp{���E�������{�=��R�;�w8O�&��=�&?����T`��u��a�E����ۖ�:�~���(5�tO���qW�{��>ٍ.���p_m�]��c���]��cQ�+��a ꓬ��6�p�APߖť�Q7�{������du�ABs��>_��<H��ܥ ���E���Ҡ����ԗpQ�#P�\{O2Z��u��0�{������]ܭ��0��hѥ���R X��eԗ���_���f�pI���a����O~�N=5�~;5�~?5�~�85�~�<5�~�:5�~�>5�~�95�~�=5�^mf�������?��ڟ�L��mf����6SB�sB�9��I�ͤ����fVhZh3-�?/��֟�̋��a.}|\g�2-�]�����n��y:���3f�S ���<#E�d�"̤�(�������g��L�b넲U��֏eu�SCã��Ⱦ>}�|�S��W�݇rؔu*�����?���<�������{��o].~I��o_���������p?=��}�a����J�J��T��<m�����}�ϛ}Y,���O��U����~L�K�I�w�#H⿼�{�6;7��WZ^��R���p3���qX0^dR�h)I�ɓ�0��2�����o����n�cP�{���7n�ң`�b�ѯD����i9_'\�P�Œ)�v�����M������t�46ԃ�Pʂ}D�ϹA�?���S2BB-T�1��@j�RH�_����n&Z=��MS���C�hZd��jt�K�`T���PJ�}:K�� e���vM���i31$�g`횖��5-���-o�������s���Tۉ��9=�Ո���;r���5���.��kD�V҅�֜���K�f[H%�IS�T�.�<UZ'R��C��.xU��L�9�ee�*t�R�Z���]*����O���JhF^��^1��GZ��R3���_%�d	q&�kJO�!��cf���	)��t��s�FmdKm�R�0 pr�[C��rŴU���(�����_�/�+���6T�ܵ�~�F�i�;f��$�A���Z����p��g��7OǕ�s��[̀qz���v{��c;����)$o�ڣ`5*�izB\>�E�5������q.�'%ŗt�0q�[�r#^�J󄧕M��EbJƝ�e�ԧshw#�N����C߳�z%�¶w����^cQ��\
n��S�a2�GhYL�`�O�
��4��9��-����L�T��fY��rl���"��ƀi~���"��ϛß��Ͼ�{��V�i�cw`<b�/�uh�3���(��f��2��9�nYRQ%��k*�p��2'��)��,tѼ����������9�.(+�Q'U�}/}w�ԗ��- VP�.�+ťla�U&�9��D��� �Y"3aܢz��X �F�h6g�W�w��|G_]���4���볯�떛�D׹��p7�_D����b���B�0�ܒ�,\8������L�<7���*�$�bt	�&��pn�w
�?��FZ)]���@���xp~sހ�gg�
Ѝ3`��v�C�﨓	-��\KK��LT�0�ŌR�bt��f�km�1�t�E���[�S&�ۓq9��X`�.�BL��f��~��gIN&���n�����_%_�e�����o0�f�K�P7`Ċ*��"OCW�h��;��u�S�	��VTI����9�E����(r��-��*�#�ZwxG�g�����FDl�u
���<�	��8$��m\P�k`���'D�V��t��!+�	��D���[�`�洠�S����I�*�*RZ�է�-L�� A.7ޯh���c�k�ʡ�?!D�9��H����T:�%F5�������y۟r���; Џ����� *��1j�h�w�V�[���P�/d�d��;�p��"UB��z- ܿ���^>R  ���N�]�B�?C�%��y��$��}��󶨁sعI^����C#'[})��M:%���^�O,�w��?�O��ߕu�������)V���n������4Wߜ/ݼڗ��o?mʏ�r��{>�Y�_�|�xx�����o�7X���j������.�����b����f�O?�S4�������l��û�ק7o�,���W���z�>��>���=ھ3�֗h���!"��l>U����7��KX�j�@�����a1C4 ,fH7���*����)2L&[�J־��B־I&S]�P��T~����B�9�����9�����=�h��
Q��Ua@�[ q���7��/�	�4h��	tԌ����yP�����Bcr��(j�fD�Z.ؙ�ͥ�Ĭ\H(���ы���D��xr�.0��V�+�Z?��F�`�!�l=ֺ��ݺdF����Y[+�Ȕ�}�L֋%"@��xz���6C�Xz�]��%��:-��0�Nd�U��pt>Q@�o6���X7�����\���l�uT������6��8H�Z���m���Bv�uwJ�,!��6&d���Y�"��$\,Ԟ䛭g[>�Z���m�)HϷ��]\��o�iT��� ���.@��]�f m�@�p:�K���Ԝ	��3�21����\�Q�ц��F�ŵ��J3j@��C2j��E��qt�k�sȀp�5�BD������������i�Y(�lf��B(jU�A�����h/*�"���xv�pѠv]D�.�C�M�䰅�$E@T!�
>�T`���LF���5j".�h�X4�6���!�lk5UD��c(j�D0��^B콇p�������	�-d�VbN6��I�M UM��`��G����" w�zFQ�3��y!���r\N��0T�\WV��V���8�!k�=q2�=�a������GOG�82�!Z,yݑYWG���Hv�	�w��'� �sE�H��[=t]�ur�N{�^E��*�1��'�`�`/ ��c88f� ��f���c7;| ��TZ�.��� ��'��c��wWcj������@�a�Ę��1B�N��j_�ԝ�D�tU9a�Wv�S=36C�X��:�uTϹ�eH�j��p�!v�$U ��C���!�;{�G�3�1�J�a+�m�(*�:[9�Ls����P����z�hc��1�g@�}� ���ź�}��d��c��e{m���Y7���J4 ��v� ��]��-(��xUf��0d�`�f����!�.����u�c��a@���X�"F�._~Au��d(U� d����C�Ga�-��|�l�@}]��ꗷ��N5���GU���s�
A��vq(�U�Eʡ�}l�Gmf�. �3��]��.��A6��:d�Lw�^ %������t�a�/����'��^�眾z������x0�b�[ ��r� �D^�Xe�����t+�k^�78�:C��'x]?! �e b#�*:���R� ~)�K�c�xwH #�@گCRW��H�1�RcW)�Y啰� �P�* �3D��r������s�:�x[DR�"J����e	 �����!�Xg�a��������';pe5��:.�s���(�69�����}u�=�L�a\��7'�m S9�
\�Zi�0�Pe�l�6�Uu*����bT��Q�W]AT��>tN�`D�:�n] �,䄴?�&����]���f��W]���p�
 i_���D듙P��i�O�������P�7��������e��>�>�����w(�?�G~�y���PK
   ���W��1W  �                  cirkitFile.jsonPK      =   �    